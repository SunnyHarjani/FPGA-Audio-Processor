-- DE1_SoC_QSYS.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DE1_SoC_QSYS is
	port (
		clk_clk                        : in    std_logic                     := '0';             --                     clk.clk
		clk_sdram_clk                  : out   std_logic;                                        --               clk_sdram.clk
		data_in_export                 : in    std_logic_vector(15 downto 0) := (others => '0'); --                 data_in.export
		data_out_export                : out   std_logic_vector(15 downto 0);                    --                data_out.export
		key_external_connection_export : in    std_logic_vector(3 downto 0)  := (others => '0'); -- key_external_connection.export
		play_btn_in_export             : in    std_logic                     := '0';             --             play_btn_in.export
		pll_locked_export              : out   std_logic;                                        --              pll_locked.export
		record_btn_in_export           : in    std_logic                     := '0';             --           record_btn_in.export
		reset_reset_n                  : in    std_logic                     := '0';             --                   reset.reset_n
		sdram_wire_addr                : out   std_logic_vector(12 downto 0);                    --              sdram_wire.addr
		sdram_wire_ba                  : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_wire_cas_n               : out   std_logic;                                        --                        .cas_n
		sdram_wire_cke                 : out   std_logic;                                        --                        .cke
		sdram_wire_cs_n                : out   std_logic;                                        --                        .cs_n
		sdram_wire_dq                  : inout std_logic_vector(15 downto 0) := (others => '0'); --                        .dq
		sdram_wire_dqm                 : out   std_logic_vector(1 downto 0);                     --                        .dqm
		sdram_wire_ras_n               : out   std_logic;                                        --                        .ras_n
		sdram_wire_we_n                : out   std_logic;                                        --                        .we_n
		sync_in_export                 : in    std_logic                     := '0'              --                 sync_in.export
	);
end entity DE1_SoC_QSYS;

architecture rtl of DE1_SoC_QSYS is
	component DE1_SoC_QSYS_PLAY_BTN_IN is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_PLAY_BTN_IN;

	component DE1_SoC_QSYS_data_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(15 downto 0) := (others => 'X')  -- export
		);
	end component DE1_SoC_QSYS_data_in;

	component DE1_SoC_QSYS_data_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component DE1_SoC_QSYS_data_out;

	component DE1_SoC_QSYS_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_jtag_uart;

	component DE1_SoC_QSYS_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_key;

	component DE1_SoC_QSYS_nios2_qsys is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(26 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component DE1_SoC_QSYS_nios2_qsys;

	component DE1_SoC_QSYS_onchip_memory2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component DE1_SoC_QSYS_onchip_memory2;

	component DE1_SoC_QSYS_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component DE1_SoC_QSYS_pll;

	component DE1_SoC_QSYS_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component DE1_SoC_QSYS_sdram;

	component DE1_SoC_QSYS_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DE1_SoC_QSYS_sysid_qsys;

	component DE1_SoC_QSYS_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component DE1_SoC_QSYS_timer;

	component DE1_SoC_QSYS_mm_interconnect_0 is
		port (
			pll_outclk0_clk                                : in  std_logic                     := 'X';             -- clk
			jtag_uart_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			nios2_qsys_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_data_master_address                 : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_qsys_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_qsys_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_qsys_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_qsys_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_instruction_master_address          : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_qsys_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_qsys_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_qsys_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			data_in_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			data_in_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			data_out_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			data_out_s1_write                              : out std_logic;                                        -- write
			data_out_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			data_out_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			data_out_s1_chipselect                         : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address            : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write              : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read               : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect         : out std_logic;                                        -- chipselect
			key_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                   : out std_logic;                                        -- write
			key_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                              : out std_logic;                                        -- chipselect
			nios2_qsys_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_qsys_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_qsys_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_memory2_s1_address                      : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_s1_write                        : out std_logic;                                        -- write
			onchip_memory2_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_s1_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory2_s1_clken                        : out std_logic;                                        -- clken
			PLAY_BTN_IN_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			PLAY_BTN_IN_s1_write                           : out std_logic;                                        -- write
			PLAY_BTN_IN_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PLAY_BTN_IN_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			PLAY_BTN_IN_s1_chipselect                      : out std_logic;                                        -- chipselect
			RECORD_BTN_IN_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			RECORD_BTN_IN_s1_write                         : out std_logic;                                        -- write
			RECORD_BTN_IN_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RECORD_BTN_IN_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			RECORD_BTN_IN_s1_chipselect                    : out std_logic;                                        -- chipselect
			sdram_s1_address                               : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                 : out std_logic;                                        -- write
			sdram_s1_read                                  : out std_logic;                                        -- read
			sdram_s1_readdata                              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                             : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                            : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                         : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                            : out std_logic;                                        -- chipselect
			sync_in_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			sync_in_s1_write                               : out std_logic;                                        -- write
			sync_in_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sync_in_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			sync_in_s1_chipselect                          : out std_logic;                                        -- chipselect
			sysid_qsys_control_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                               : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                                 : out std_logic;                                        -- write
			timer_s1_readdata                              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                             : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                            : out std_logic                                         -- chipselect
		);
	end component DE1_SoC_QSYS_mm_interconnect_0;

	component DE1_SoC_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component DE1_SoC_QSYS_irq_mapper;

	component de1_soc_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component de1_soc_qsys_rst_controller;

	component de1_soc_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component de1_soc_qsys_rst_controller_001;

	signal pll_outclk0_clk                                               : std_logic;                     -- pll:outclk_0 -> [PLAY_BTN_IN:clk, RECORD_BTN_IN:clk, data_in:clk, data_out:clk, irq_mapper:clk, jtag_uart:clk, key:clk, mm_interconnect_0:pll_outclk0_clk, nios2_qsys:clk, onchip_memory2:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sync_in:clk, sysid_qsys:clock, timer:clk]
	signal nios2_qsys_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	signal nios2_qsys_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	signal nios2_qsys_data_master_debugaccess                            : std_logic;                     -- nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	signal nios2_qsys_data_master_address                                : std_logic_vector(26 downto 0); -- nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	signal nios2_qsys_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	signal nios2_qsys_data_master_read                                   : std_logic;                     -- nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	signal nios2_qsys_data_master_write                                  : std_logic;                     -- nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	signal nios2_qsys_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	signal nios2_qsys_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	signal nios2_qsys_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	signal nios2_qsys_instruction_master_address                         : std_logic_vector(26 downto 0); -- nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	signal nios2_qsys_instruction_master_read                            : std_logic;                     -- nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_qsys_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata       : std_logic_vector(31 downto 0); -- nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest    : std_logic;                     -- nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess    : std_logic;                     -- mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_address        : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_read           : std_logic;                     -- mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_write          : std_logic;                     -- mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	signal mm_interconnect_0_onchip_memory2_s1_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	signal mm_interconnect_0_onchip_memory2_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	signal mm_interconnect_0_onchip_memory2_s1_address                   : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	signal mm_interconnect_0_onchip_memory2_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	signal mm_interconnect_0_onchip_memory2_s1_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	signal mm_interconnect_0_onchip_memory2_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	signal mm_interconnect_0_onchip_memory2_s1_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	signal mm_interconnect_0_timer_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                           : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_0:timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_s1_address -> timer:address
	signal mm_interconnect_0_timer_s1_write                              : std_logic;                     -- mm_interconnect_0:timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_0_key_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_readdata                             : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_write                                : std_logic;                     -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                           : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                        : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                            : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                               : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                      : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                              : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_sync_in_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:sync_in_s1_chipselect -> sync_in:chipselect
	signal mm_interconnect_0_sync_in_s1_readdata                         : std_logic_vector(31 downto 0); -- sync_in:readdata -> mm_interconnect_0:sync_in_s1_readdata
	signal mm_interconnect_0_sync_in_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sync_in_s1_address -> sync_in:address
	signal mm_interconnect_0_sync_in_s1_write                            : std_logic;                     -- mm_interconnect_0:sync_in_s1_write -> mm_interconnect_0_sync_in_s1_write:in
	signal mm_interconnect_0_sync_in_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sync_in_s1_writedata -> sync_in:writedata
	signal mm_interconnect_0_data_out_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:data_out_s1_chipselect -> data_out:chipselect
	signal mm_interconnect_0_data_out_s1_readdata                        : std_logic_vector(31 downto 0); -- data_out:readdata -> mm_interconnect_0:data_out_s1_readdata
	signal mm_interconnect_0_data_out_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:data_out_s1_address -> data_out:address
	signal mm_interconnect_0_data_out_s1_write                           : std_logic;                     -- mm_interconnect_0:data_out_s1_write -> mm_interconnect_0_data_out_s1_write:in
	signal mm_interconnect_0_data_out_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:data_out_s1_writedata -> data_out:writedata
	signal mm_interconnect_0_data_in_s1_readdata                         : std_logic_vector(31 downto 0); -- data_in:readdata -> mm_interconnect_0:data_in_s1_readdata
	signal mm_interconnect_0_data_in_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:data_in_s1_address -> data_in:address
	signal mm_interconnect_0_play_btn_in_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:PLAY_BTN_IN_s1_chipselect -> PLAY_BTN_IN:chipselect
	signal mm_interconnect_0_play_btn_in_s1_readdata                     : std_logic_vector(31 downto 0); -- PLAY_BTN_IN:readdata -> mm_interconnect_0:PLAY_BTN_IN_s1_readdata
	signal mm_interconnect_0_play_btn_in_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PLAY_BTN_IN_s1_address -> PLAY_BTN_IN:address
	signal mm_interconnect_0_play_btn_in_s1_write                        : std_logic;                     -- mm_interconnect_0:PLAY_BTN_IN_s1_write -> mm_interconnect_0_play_btn_in_s1_write:in
	signal mm_interconnect_0_play_btn_in_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:PLAY_BTN_IN_s1_writedata -> PLAY_BTN_IN:writedata
	signal mm_interconnect_0_record_btn_in_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:RECORD_BTN_IN_s1_chipselect -> RECORD_BTN_IN:chipselect
	signal mm_interconnect_0_record_btn_in_s1_readdata                   : std_logic_vector(31 downto 0); -- RECORD_BTN_IN:readdata -> mm_interconnect_0:RECORD_BTN_IN_s1_readdata
	signal mm_interconnect_0_record_btn_in_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:RECORD_BTN_IN_s1_address -> RECORD_BTN_IN:address
	signal mm_interconnect_0_record_btn_in_s1_write                      : std_logic;                     -- mm_interconnect_0:RECORD_BTN_IN_s1_write -> mm_interconnect_0_record_btn_in_s1_write:in
	signal mm_interconnect_0_record_btn_in_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:RECORD_BTN_IN_s1_writedata -> RECORD_BTN_IN:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- timer:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- key:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- sync_in:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                      : std_logic;                     -- PLAY_BTN_IN:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                      : std_logic;                     -- RECORD_BTN_IN:irq -> irq_mapper:receiver5_irq
	signal nios2_qsys_d_irq_irq                                          : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys:d_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                        : std_logic;                     -- rst_controller_001:reset_req -> [nios2_qsys:reset_req, rst_translator_001:reset_req_in]
	signal nios2_qsys_jtag_debug_module_reset_reset                      : std_logic;                     -- nios2_qsys:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [pll:rst, rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                     : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv               : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_sync_in_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_sync_in_s1_write:inv -> sync_in:write_n
	signal mm_interconnect_0_data_out_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_data_out_s1_write:inv -> data_out:write_n
	signal mm_interconnect_0_play_btn_in_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_play_btn_in_s1_write:inv -> PLAY_BTN_IN:write_n
	signal mm_interconnect_0_record_btn_in_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_record_btn_in_s1_write:inv -> RECORD_BTN_IN:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [PLAY_BTN_IN:reset_n, RECORD_BTN_IN:reset_n, data_in:reset_n, data_out:reset_n, jtag_uart:rst_n, key:reset_n, sdram:reset_n, sync_in:reset_n, sysid_qsys:reset_n, timer:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> nios2_qsys:reset_n

begin

	play_btn_in : component DE1_SoC_QSYS_PLAY_BTN_IN
		port map (
			clk        => pll_outclk0_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_play_btn_in_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_play_btn_in_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_play_btn_in_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_play_btn_in_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_play_btn_in_s1_readdata,        --                    .readdata
			in_port    => play_btn_in_export,                               -- external_connection.export
			irq        => irq_mapper_receiver4_irq                          --                 irq.irq
		);

	record_btn_in : component DE1_SoC_QSYS_PLAY_BTN_IN
		port map (
			clk        => pll_outclk0_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_record_btn_in_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_record_btn_in_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_record_btn_in_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_record_btn_in_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_record_btn_in_s1_readdata,        --                    .readdata
			in_port    => record_btn_in_export,                               -- external_connection.export
			irq        => irq_mapper_receiver5_irq                            --                 irq.irq
		);

	data_in : component DE1_SoC_QSYS_data_in
		port map (
			clk      => pll_outclk0_clk,                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_data_in_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_data_in_s1_readdata,    --                    .readdata
			in_port  => data_in_export                            -- external_connection.export
		);

	data_out : component DE1_SoC_QSYS_data_out
		port map (
			clk        => pll_outclk0_clk,                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_data_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_data_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_data_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_data_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_data_out_s1_readdata,        --                    .readdata
			out_port   => data_out_export                                -- external_connection.export
		);

	jtag_uart : component DE1_SoC_QSYS_jtag_uart
		port map (
			clk            => pll_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	key : component DE1_SoC_QSYS_key
		port map (
			clk        => pll_outclk0_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port    => key_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                  --                 irq.irq
		);

	nios2_qsys : component DE1_SoC_QSYS_nios2_qsys
		port map (
			clk                                   => pll_outclk0_clk,                                            --                       clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,               --                   reset_n.reset_n
			reset_req                             => rst_controller_001_reset_out_reset_req,                     --                          .reset_req
			d_address                             => nios2_qsys_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_qsys_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2 : component DE1_SoC_QSYS_onchip_memory2
		port map (
			clk        => pll_outclk0_clk,                                --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,             --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	pll : component DE1_SoC_QSYS_pll
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_outclk0_clk,         -- outclk0.clk
			outclk_1 => clk_sdram_clk,           -- outclk1.clk
			locked   => pll_locked_export        --  locked.export
		);

	sdram : component DE1_SoC_QSYS_sdram
		port map (
			clk            => pll_outclk0_clk,                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	sync_in : component DE1_SoC_QSYS_PLAY_BTN_IN
		port map (
			clk        => pll_outclk0_clk,                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_sync_in_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sync_in_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sync_in_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sync_in_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sync_in_s1_readdata,        --                    .readdata
			in_port    => sync_in_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                      --                 irq.irq
		);

	sysid_qsys : component DE1_SoC_QSYS_sysid_qsys
		port map (
			clock    => pll_outclk0_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_control_slave_address(0)  --              .address
		);

	timer : component DE1_SoC_QSYS_timer
		port map (
			clk        => pll_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                    --   irq.irq
		);

	mm_interconnect_0 : component DE1_SoC_QSYS_mm_interconnect_0
		port map (
			pll_outclk0_clk                                => pll_outclk0_clk,                                            --                              pll_outclk0.clk
			jtag_uart_reset_reset_bridge_in_reset_reset    => rst_controller_reset_out_reset,                             --    jtag_uart_reset_reset_bridge_in_reset.reset
			nios2_qsys_reset_n_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                         -- nios2_qsys_reset_n_reset_bridge_in_reset.reset
			nios2_qsys_data_master_address                 => nios2_qsys_data_master_address,                             --                   nios2_qsys_data_master.address
			nios2_qsys_data_master_waitrequest             => nios2_qsys_data_master_waitrequest,                         --                                         .waitrequest
			nios2_qsys_data_master_byteenable              => nios2_qsys_data_master_byteenable,                          --                                         .byteenable
			nios2_qsys_data_master_read                    => nios2_qsys_data_master_read,                                --                                         .read
			nios2_qsys_data_master_readdata                => nios2_qsys_data_master_readdata,                            --                                         .readdata
			nios2_qsys_data_master_write                   => nios2_qsys_data_master_write,                               --                                         .write
			nios2_qsys_data_master_writedata               => nios2_qsys_data_master_writedata,                           --                                         .writedata
			nios2_qsys_data_master_debugaccess             => nios2_qsys_data_master_debugaccess,                         --                                         .debugaccess
			nios2_qsys_instruction_master_address          => nios2_qsys_instruction_master_address,                      --            nios2_qsys_instruction_master.address
			nios2_qsys_instruction_master_waitrequest      => nios2_qsys_instruction_master_waitrequest,                  --                                         .waitrequest
			nios2_qsys_instruction_master_read             => nios2_qsys_instruction_master_read,                         --                                         .read
			nios2_qsys_instruction_master_readdata         => nios2_qsys_instruction_master_readdata,                     --                                         .readdata
			data_in_s1_address                             => mm_interconnect_0_data_in_s1_address,                       --                               data_in_s1.address
			data_in_s1_readdata                            => mm_interconnect_0_data_in_s1_readdata,                      --                                         .readdata
			data_out_s1_address                            => mm_interconnect_0_data_out_s1_address,                      --                              data_out_s1.address
			data_out_s1_write                              => mm_interconnect_0_data_out_s1_write,                        --                                         .write
			data_out_s1_readdata                           => mm_interconnect_0_data_out_s1_readdata,                     --                                         .readdata
			data_out_s1_writedata                          => mm_interconnect_0_data_out_s1_writedata,                    --                                         .writedata
			data_out_s1_chipselect                         => mm_interconnect_0_data_out_s1_chipselect,                   --                                         .chipselect
			jtag_uart_avalon_jtag_slave_address            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,      --              jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,        --                                         .write
			jtag_uart_avalon_jtag_slave_read               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,         --                                         .read
			jtag_uart_avalon_jtag_slave_readdata           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,     --                                         .readdata
			jtag_uart_avalon_jtag_slave_writedata          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,    --                                         .writedata
			jtag_uart_avalon_jtag_slave_waitrequest        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,  --                                         .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,   --                                         .chipselect
			key_s1_address                                 => mm_interconnect_0_key_s1_address,                           --                                   key_s1.address
			key_s1_write                                   => mm_interconnect_0_key_s1_write,                             --                                         .write
			key_s1_readdata                                => mm_interconnect_0_key_s1_readdata,                          --                                         .readdata
			key_s1_writedata                               => mm_interconnect_0_key_s1_writedata,                         --                                         .writedata
			key_s1_chipselect                              => mm_interconnect_0_key_s1_chipselect,                        --                                         .chipselect
			nios2_qsys_jtag_debug_module_address           => mm_interconnect_0_nios2_qsys_jtag_debug_module_address,     --             nios2_qsys_jtag_debug_module.address
			nios2_qsys_jtag_debug_module_write             => mm_interconnect_0_nios2_qsys_jtag_debug_module_write,       --                                         .write
			nios2_qsys_jtag_debug_module_read              => mm_interconnect_0_nios2_qsys_jtag_debug_module_read,        --                                         .read
			nios2_qsys_jtag_debug_module_readdata          => mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata,    --                                         .readdata
			nios2_qsys_jtag_debug_module_writedata         => mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata,   --                                         .writedata
			nios2_qsys_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable,  --                                         .byteenable
			nios2_qsys_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest, --                                         .waitrequest
			nios2_qsys_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess, --                                         .debugaccess
			onchip_memory2_s1_address                      => mm_interconnect_0_onchip_memory2_s1_address,                --                        onchip_memory2_s1.address
			onchip_memory2_s1_write                        => mm_interconnect_0_onchip_memory2_s1_write,                  --                                         .write
			onchip_memory2_s1_readdata                     => mm_interconnect_0_onchip_memory2_s1_readdata,               --                                         .readdata
			onchip_memory2_s1_writedata                    => mm_interconnect_0_onchip_memory2_s1_writedata,              --                                         .writedata
			onchip_memory2_s1_byteenable                   => mm_interconnect_0_onchip_memory2_s1_byteenable,             --                                         .byteenable
			onchip_memory2_s1_chipselect                   => mm_interconnect_0_onchip_memory2_s1_chipselect,             --                                         .chipselect
			onchip_memory2_s1_clken                        => mm_interconnect_0_onchip_memory2_s1_clken,                  --                                         .clken
			PLAY_BTN_IN_s1_address                         => mm_interconnect_0_play_btn_in_s1_address,                   --                           PLAY_BTN_IN_s1.address
			PLAY_BTN_IN_s1_write                           => mm_interconnect_0_play_btn_in_s1_write,                     --                                         .write
			PLAY_BTN_IN_s1_readdata                        => mm_interconnect_0_play_btn_in_s1_readdata,                  --                                         .readdata
			PLAY_BTN_IN_s1_writedata                       => mm_interconnect_0_play_btn_in_s1_writedata,                 --                                         .writedata
			PLAY_BTN_IN_s1_chipselect                      => mm_interconnect_0_play_btn_in_s1_chipselect,                --                                         .chipselect
			RECORD_BTN_IN_s1_address                       => mm_interconnect_0_record_btn_in_s1_address,                 --                         RECORD_BTN_IN_s1.address
			RECORD_BTN_IN_s1_write                         => mm_interconnect_0_record_btn_in_s1_write,                   --                                         .write
			RECORD_BTN_IN_s1_readdata                      => mm_interconnect_0_record_btn_in_s1_readdata,                --                                         .readdata
			RECORD_BTN_IN_s1_writedata                     => mm_interconnect_0_record_btn_in_s1_writedata,               --                                         .writedata
			RECORD_BTN_IN_s1_chipselect                    => mm_interconnect_0_record_btn_in_s1_chipselect,              --                                         .chipselect
			sdram_s1_address                               => mm_interconnect_0_sdram_s1_address,                         --                                 sdram_s1.address
			sdram_s1_write                                 => mm_interconnect_0_sdram_s1_write,                           --                                         .write
			sdram_s1_read                                  => mm_interconnect_0_sdram_s1_read,                            --                                         .read
			sdram_s1_readdata                              => mm_interconnect_0_sdram_s1_readdata,                        --                                         .readdata
			sdram_s1_writedata                             => mm_interconnect_0_sdram_s1_writedata,                       --                                         .writedata
			sdram_s1_byteenable                            => mm_interconnect_0_sdram_s1_byteenable,                      --                                         .byteenable
			sdram_s1_readdatavalid                         => mm_interconnect_0_sdram_s1_readdatavalid,                   --                                         .readdatavalid
			sdram_s1_waitrequest                           => mm_interconnect_0_sdram_s1_waitrequest,                     --                                         .waitrequest
			sdram_s1_chipselect                            => mm_interconnect_0_sdram_s1_chipselect,                      --                                         .chipselect
			sync_in_s1_address                             => mm_interconnect_0_sync_in_s1_address,                       --                               sync_in_s1.address
			sync_in_s1_write                               => mm_interconnect_0_sync_in_s1_write,                         --                                         .write
			sync_in_s1_readdata                            => mm_interconnect_0_sync_in_s1_readdata,                      --                                         .readdata
			sync_in_s1_writedata                           => mm_interconnect_0_sync_in_s1_writedata,                     --                                         .writedata
			sync_in_s1_chipselect                          => mm_interconnect_0_sync_in_s1_chipselect,                    --                                         .chipselect
			sysid_qsys_control_slave_address               => mm_interconnect_0_sysid_qsys_control_slave_address,         --                 sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata              => mm_interconnect_0_sysid_qsys_control_slave_readdata,        --                                         .readdata
			timer_s1_address                               => mm_interconnect_0_timer_s1_address,                         --                                 timer_s1.address
			timer_s1_write                                 => mm_interconnect_0_timer_s1_write,                           --                                         .write
			timer_s1_readdata                              => mm_interconnect_0_timer_s1_readdata,                        --                                         .readdata
			timer_s1_writedata                             => mm_interconnect_0_timer_s1_writedata,                       --                                         .writedata
			timer_s1_chipselect                            => mm_interconnect_0_timer_s1_chipselect                       --                                         .chipselect
		);

	irq_mapper : component DE1_SoC_QSYS_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                    --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			sender_irq    => nios2_qsys_d_irq_irq                --    sender.irq
		);

	rst_controller : component de1_soc_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_outclk0_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component de1_soc_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                  -- reset_in0.reset
			reset_in1      => nios2_qsys_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => pll_outclk0_clk,                          --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_sync_in_s1_write_ports_inv <= not mm_interconnect_0_sync_in_s1_write;

	mm_interconnect_0_data_out_s1_write_ports_inv <= not mm_interconnect_0_data_out_s1_write;

	mm_interconnect_0_play_btn_in_s1_write_ports_inv <= not mm_interconnect_0_play_btn_in_s1_write;

	mm_interconnect_0_record_btn_in_s1_write_ports_inv <= not mm_interconnect_0_record_btn_in_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of DE1_SoC_QSYS
